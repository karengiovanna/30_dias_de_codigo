LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY P_xor IS
  PORT(
    in_port_A : IN STD_LOGIC;
    in_port_B : IN STD_LOGIC;
    out_port  : OUT STD_LOGIC
    );
END ENTITY;
